//cpu, descricao da controle operativo

module NRISC_CPU(
				
				)
endmodule;