//ULA


module NRISC_ULA(
					ULA_A, //ULA input A
					ULA_B, //ULA input B
					ULA_OUT,
					ULA_ctrl,
					ULA_flags,
					clk,
					rst					
					);

endmodule;